module pseudo_random_gen
(
  // Clock and Reset
  input  logic        clk,
  input  logic        rst,

  output wire        fault,
  output wire        index
);

endmodule
